----
-- @author: Douglas Martins, Lucas M. Mendes, Matheus R. Willemann
-- Projeto Final ELD - gerador de Figuras de Lissajous

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

--library ieee_proposed;
--use iee_proposed.fixed_pkg.all;


--- TODO: ver lookup table funções Sin e cos ou implementação polinomial

entity lissajous_curves is
  port(
    x_out, y_out  : out std_logic_vector(15 downto 0) := X"0000" ; -- inteiros de 16 bits
    var_in : in std_logic_vector(15 downto 0);
    next_bt : in std_logic;
    clk: in std_logic
);
end lissajous_curves;

-- Este sistema utiliza um sistema numérico de ponto fixo, com número de casas
-- decimais dado por dec_offset

  --TODO: fazer process para ajustar valores das variaveis

architecture arq of lissajous_curves is

  -- tipos
-- constant precision : integer := 32;
  subtype int is signed(31 downto 0);

  -- Constantes
  constant pi : integer := 3141; -- pi with decimal offset
  constant dec_offset : integer := 1000;

  -- Variáveis
  shared variable x_ampl  : integer := 5000; -- 5v
  shared variable y_ampl  : integer := 5000;
  shared variable alpha   : integer := 2000;
  shared variable beta    : integer := 4000;
  shared variable delta   : integer := 0;
  shared variable t       : integer := 0;
	shared variable x_tmp   : std_logic_vector(15 downto 0);
	shared variable y_tmp   : std_logic_vector(15 downto 0);

-- Funções

  -- Multiplicação, levando em conta o offset decimal
  pure function mult (x: integer; y : integer) return integer is
  begin
    return (x*y)/dec_offset;
  end function;
  -- Divisao
  pure function div (x: integer; y : integer) return integer is
  begin
    return (x*dec_offset)/y;
  end function;

  -- Aproximação de Taylor de seno, com boa precisão entre 0 e 90º
--   pure function sin_0_pi2 (x : int) return int is
--     constant t_3 : int := to_signed(6,32)*dec_offset; -- 6*dec_offset;
--     constant t_5 : int := to_signed(120,32)*dec_offset;-- 120*dec_offset;
--   begin
--     return x - div( mult(x,mult(x,x)) , t_3) + div( mult(x,mult(x,mult(x,mult(x,x)))), t_5);
--   end function;

--   pure function sin (x : int := "0") return int is
--     variable quadrant :  int := "00";
--     --variable angl : integer := angle mod 360;
-- begin

--   quadrant := div(x, pi/2);
--   case quadrant is
--     when "00" =>
--       return sin_0_pi2(x);
--     when "01" =>
--       return sin_0_pi2(x-pi);
--     when "10" =>
--       return -1*sin_0_pi2(x);
--     when others =>
--       return -1*sin_0_pi2(x-pi);
--   end case;
-- end function;

  -- Seno implementado por tabela
  function sin_0_pi2 ( rad : integer ) return integer is
  begin
    case rad is
      when  0  => return  0 ;
      when  1  => return  1 ;
      when  2  => return  2 ;
      when  3  => return  3 ;
      when  4  => return  4 ;
      when  5  => return  5 ;
      when  6  => return  6 ;
      when  7  => return  7 ;
      when  8  => return  8 ;
      when  9  => return  9 ;
      when  10  => return  10 ;
      when  11  => return  11 ;
      when  12  => return  12 ;
      when  13  => return  13 ;
      when  14  => return  14 ;
      when  15  => return  15 ;
      when  16  => return  16 ;
      when  17  => return  17 ;
      when  18  => return  18 ;
      when  19  => return  19 ;
      when  20  => return  20 ;
      when  21  => return  21 ;
      when  22  => return  22 ;
      when  23  => return  23 ;
      when  24  => return  24 ;
      when  25  => return  25 ;
      when  26  => return  26 ;
      when  27  => return  27 ;
      when  28  => return  28 ;
      when  29  => return  29 ;
      when  30  => return  30 ;
      when  31  => return  31 ;
      when  32  => return  32 ;
      when  33  => return  33 ;
      when  34  => return  34 ;
      when  35  => return  35 ;
      when  36  => return  36 ;
      when  37  => return  37 ;
      when  38  => return  38 ;
      when  39  => return  39 ;
      when  40  => return  40 ;
      when  41  => return  41 ;
      when  42  => return  42 ;
      when  43  => return  43 ;
      when  44  => return  44 ;
      when  45  => return  45 ;
      when  46  => return  46 ;
      when  47  => return  47 ;
      when  48  => return  48 ;
      when  49  => return  49 ;
      when  50  => return  50 ;
      when  51  => return  51 ;
      when  52  => return  52 ;
      when  53  => return  53 ;
      when  54  => return  54 ;
      when  55  => return  55 ;
      when  56  => return  56 ;
      when  57  => return  57 ;
      when  58  => return  58 ;
      when  59  => return  59 ;
      when  60  => return  60 ;
      when  61  => return  61 ;
      when  62  => return  62 ;
      when  63  => return  63 ;
      when  64  => return  64 ;
      when  65  => return  65 ;
      when  66  => return  66 ;
      when  67  => return  67 ;
      when  68  => return  68 ;
      when  69  => return  69 ;
      when  70  => return  70 ;
      when  71  => return  71 ;
      when  72  => return  72 ;
      when  73  => return  73 ;
      when  74  => return  74 ;
      when  75  => return  75 ;
      when  76  => return  76 ;
      when  77  => return  77 ;
      when  78  => return  78 ;
      when  79  => return  79 ;
      when  80  => return  80 ;
      when  81  => return  81 ;
      when  82  => return  82 ;
      when  83  => return  83 ;
      when  84  => return  84 ;
      when  85  => return  85 ;
      when  86  => return  86 ;
      when  87  => return  87 ;
      when  88  => return  88 ;
      when  89  => return  89 ;
      when  90  => return  90 ;
      when  91  => return  91 ;
      when  92  => return  92 ;
      when  93  => return  93 ;
      when  94  => return  94 ;
      when  95  => return  95 ;
      when  96  => return  96 ;
      when  97  => return  97 ;
      when  98  => return  98 ;
      when  99  => return  99 ;
      when  100  => return  100 ;
      when  101  => return  101 ;
      when  102  => return  102 ;
      when  103  => return  103 ;
      when  104  => return  104 ;
      when  105  => return  105 ;
      when  106  => return  106 ;
      when  107  => return  107 ;
      when  108  => return  108 ;
      when  109  => return  109 ;
      when  110  => return  110 ;
      when  111  => return  111 ;
      when  112  => return  112 ;
      when  113  => return  113 ;
      when  114  => return  114 ;
      when  115  => return  115 ;
      when  116  => return  116 ;
      when  117  => return  117 ;
      when  118  => return  118 ;
      when  119  => return  119 ;
      when  120  => return  120 ;
      when  121  => return  121 ;
      when  122  => return  122 ;
      when  123  => return  123 ;
      when  124  => return  124 ;
      when  125  => return  125 ;
      when  126  => return  126 ;
      when  127  => return  127 ;
      when  128  => return  128 ;
      when  129  => return  129 ;
      when  130  => return  130 ;
      when  131  => return  131 ;
      when  132  => return  132 ;
      when  133  => return  133 ;
      when  134  => return  134 ;
      when  135  => return  135 ;
      when  136  => return  136 ;
      when  137  => return  137 ;
      when  138  => return  138 ;
      when  139  => return  139 ;
      when  140  => return  140 ;
      when  141  => return  141 ;
      when  142  => return  142 ;
      when  143  => return  143 ;
      when  144  => return  144 ;
      when  145  => return  144 ;
      when  146  => return  145 ;
      when  147  => return  146 ;
      when  148  => return  147 ;
      when  149  => return  148 ;
      when  150  => return  149 ;
      when  151  => return  150 ;
      when  152  => return  151 ;
      when  153  => return  152 ;
      when  154  => return  153 ;
      when  155  => return  154 ;
      when  156  => return  155 ;
      when  157  => return  156 ;
      when  158  => return  157 ;
      when  159  => return  158 ;
      when  160  => return  159 ;
      when  161  => return  160 ;
      when  162  => return  161 ;
      when  163  => return  162 ;
      when  164  => return  163 ;
      when  165  => return  164 ;
      when  166  => return  165 ;
      when  167  => return  166 ;
      when  168  => return  167 ;
      when  169  => return  168 ;
      when  170  => return  169 ;
      when  171  => return  170 ;
      when  172  => return  171 ;
      when  173  => return  172 ;
      when  174  => return  173 ;
      when  175  => return  174 ;
      when  176  => return  175 ;
      when  177  => return  176 ;
      when  178  => return  177 ;
      when  179  => return  178 ;
      when  180  => return  179 ;
      when  181  => return  180 ;
      when  182  => return  181 ;
      when  183  => return  182 ;
      when  184  => return  183 ;
      when  185  => return  184 ;
      when  186  => return  185 ;
      when  187  => return  186 ;
      when  188  => return  187 ;
      when  189  => return  188 ;
      when  190  => return  189 ;
      when  191  => return  190 ;
      when  192  => return  191 ;
      when  193  => return  192 ;
      when  194  => return  193 ;
      when  195  => return  194 ;
      when  196  => return  195 ;
      when  197  => return  196 ;
      when  198  => return  197 ;
      when  199  => return  198 ;
      when  200  => return  199 ;
      when  201  => return  200 ;
      when  202  => return  201 ;
      when  203  => return  202 ;
      when  204  => return  203 ;
      when  205  => return  204 ;
      when  206  => return  205 ;
      when  207  => return  206 ;
      when  208  => return  207 ;
      when  209  => return  207 ;
      when  210  => return  208 ;
      when  211  => return  209 ;
      when  212  => return  210 ;
      when  213  => return  211 ;
      when  214  => return  212 ;
      when  215  => return  213 ;
      when  216  => return  214 ;
      when  217  => return  215 ;
      when  218  => return  216 ;
      when  219  => return  217 ;
      when  220  => return  218 ;
      when  221  => return  219 ;
      when  222  => return  220 ;
      when  223  => return  221 ;
      when  224  => return  222 ;
      when  225  => return  223 ;
      when  226  => return  224 ;
      when  227  => return  225 ;
      when  228  => return  226 ;
      when  229  => return  227 ;
      when  230  => return  228 ;
      when  231  => return  229 ;
      when  232  => return  230 ;
      when  233  => return  231 ;
      when  234  => return  232 ;
      when  235  => return  233 ;
      when  236  => return  234 ;
      when  237  => return  235 ;
      when  238  => return  236 ;
      when  239  => return  237 ;
      when  240  => return  238 ;
      when  241  => return  239 ;
      when  242  => return  240 ;
      when  243  => return  241 ;
      when  244  => return  242 ;
      when  245  => return  243 ;
      when  246  => return  244 ;
      when  247  => return  244 ;
      when  248  => return  245 ;
      when  249  => return  246 ;
      when  250  => return  247 ;
      when  251  => return  248 ;
      when  252  => return  249 ;
      when  253  => return  250 ;
      when  254  => return  251 ;
      when  255  => return  252 ;
      when  256  => return  253 ;
      when  257  => return  254 ;
      when  258  => return  255 ;
      when  259  => return  256 ;
      when  260  => return  257 ;
      when  261  => return  258 ;
      when  262  => return  259 ;
      when  263  => return  260 ;
      when  264  => return  261 ;
      when  265  => return  262 ;
      when  266  => return  263 ;
      when  267  => return  264 ;
      when  268  => return  265 ;
      when  269  => return  266 ;
      when  270  => return  267 ;
      when  271  => return  268 ;
      when  272  => return  269 ;
      when  273  => return  270 ;
      when  274  => return  271 ;
      when  275  => return  272 ;
      when  276  => return  273 ;
      when  277  => return  273 ;
      when  278  => return  274 ;
      when  279  => return  275 ;
      when  280  => return  276 ;
      when  281  => return  277 ;
      when  282  => return  278 ;
      when  283  => return  279 ;
      when  284  => return  280 ;
      when  285  => return  281 ;
      when  286  => return  282 ;
      when  287  => return  283 ;
      when  288  => return  284 ;
      when  289  => return  285 ;
      when  290  => return  286 ;
      when  291  => return  287 ;
      when  292  => return  288 ;
      when  293  => return  289 ;
      when  294  => return  290 ;
      when  295  => return  291 ;
      when  296  => return  292 ;
      when  297  => return  293 ;
      when  298  => return  294 ;
      when  299  => return  295 ;
      when  300  => return  296 ;
      when  301  => return  296 ;
      when  302  => return  297 ;
      when  303  => return  298 ;
      when  304  => return  299 ;
      when  305  => return  300 ;
      when  306  => return  301 ;
      when  307  => return  302 ;
      when  308  => return  303 ;
      when  309  => return  304 ;
      when  310  => return  305 ;
      when  311  => return  306 ;
      when  312  => return  307 ;
      when  313  => return  308 ;
      when  314  => return  309 ;
      when  315  => return  310 ;
      when  316  => return  311 ;
      when  317  => return  312 ;
      when  318  => return  313 ;
      when  319  => return  314 ;
      when  320  => return  315 ;
      when  321  => return  316 ;
      when  322  => return  316 ;
      when  323  => return  317 ;
      when  324  => return  318 ;
      when  325  => return  319 ;
      when  326  => return  320 ;
      when  327  => return  321 ;
      when  328  => return  322 ;
      when  329  => return  323 ;
      when  330  => return  324 ;
      when  331  => return  325 ;
      when  332  => return  326 ;
      when  333  => return  327 ;
      when  334  => return  328 ;
      when  335  => return  329 ;
      when  336  => return  330 ;
      when  337  => return  331 ;
      when  338  => return  332 ;
      when  339  => return  333 ;
      when  340  => return  333 ;
      when  341  => return  334 ;
      when  342  => return  335 ;
      when  343  => return  336 ;
      when  344  => return  337 ;
      when  345  => return  338 ;
      when  346  => return  339 ;
      when  347  => return  340 ;
      when  348  => return  341 ;
      when  349  => return  342 ;
      when  350  => return  343 ;
      when  351  => return  344 ;
      when  352  => return  345 ;
      when  353  => return  346 ;
      when  354  => return  347 ;
      when  355  => return  348 ;
      when  356  => return  349 ;
      when  357  => return  349 ;
      when  358  => return  350 ;
      when  359  => return  351 ;
      when  360  => return  352 ;
      when  361  => return  353 ;
      when  362  => return  354 ;
      when  363  => return  355 ;
      when  364  => return  356 ;
      when  365  => return  357 ;
      when  366  => return  358 ;
      when  367  => return  359 ;
      when  368  => return  360 ;
      when  369  => return  361 ;
      when  370  => return  362 ;
      when  371  => return  363 ;
      when  372  => return  363 ;
      when  373  => return  364 ;
      when  374  => return  365 ;
      when  375  => return  366 ;
      when  376  => return  367 ;
      when  377  => return  368 ;
      when  378  => return  369 ;
      when  379  => return  370 ;
      when  380  => return  371 ;
      when  381  => return  372 ;
      when  382  => return  373 ;
      when  383  => return  374 ;
      when  384  => return  375 ;
      when  385  => return  376 ;
      when  386  => return  376 ;
      when  387  => return  377 ;
      when  388  => return  378 ;
      when  389  => return  379 ;
      when  390  => return  380 ;
      when  391  => return  381 ;
      when  392  => return  382 ;
      when  393  => return  383 ;
      when  394  => return  384 ;
      when  395  => return  385 ;
      when  396  => return  386 ;
      when  397  => return  387 ;
      when  398  => return  388 ;
      when  399  => return  388 ;
      when  400  => return  389 ;
      when  401  => return  390 ;
      when  402  => return  391 ;
      when  403  => return  392 ;
      when  404  => return  393 ;
      when  405  => return  394 ;
      when  406  => return  395 ;
      when  407  => return  396 ;
      when  408  => return  397 ;
      when  409  => return  398 ;
      when  410  => return  399 ;
      when  411  => return  400 ;
      when  412  => return  400 ;
      when  413  => return  401 ;
      when  414  => return  402 ;
      when  415  => return  403 ;
      when  416  => return  404 ;
      when  417  => return  405 ;
      when  418  => return  406 ;
      when  419  => return  407 ;
      when  420  => return  408 ;
      when  421  => return  409 ;
      when  422  => return  410 ;
      when  423  => return  410 ;
      when  424  => return  411 ;
      when  425  => return  412 ;
      when  426  => return  413 ;
      when  427  => return  414 ;
      when  428  => return  415 ;
      when  429  => return  416 ;
      when  430  => return  417 ;
      when  431  => return  418 ;
      when  432  => return  419 ;
      when  433  => return  420 ;
      when  434  => return  421 ;
      when  435  => return  421 ;
      when  436  => return  422 ;
      when  437  => return  423 ;
      when  438  => return  424 ;
      when  439  => return  425 ;
      when  440  => return  426 ;
      when  441  => return  427 ;
      when  442  => return  428 ;
      when  443  => return  429 ;
      when  444  => return  430 ;
      when  445  => return  430 ;
      when  446  => return  431 ;
      when  447  => return  432 ;
      when  448  => return  433 ;
      when  449  => return  434 ;
      when  450  => return  435 ;
      when  451  => return  436 ;
      when  452  => return  437 ;
      when  453  => return  438 ;
      when  454  => return  439 ;
      when  455  => return  439 ;
      when  456  => return  440 ;
      when  457  => return  441 ;
      when  458  => return  442 ;
      when  459  => return  443 ;
      when  460  => return  444 ;
      when  461  => return  445 ;
      when  462  => return  446 ;
      when  463  => return  447 ;
      when  464  => return  448 ;
      when  465  => return  448 ;
      when  466  => return  449 ;
      when  467  => return  450 ;
      when  468  => return  451 ;
      when  469  => return  452 ;
      when  470  => return  453 ;
      when  471  => return  454 ;
      when  472  => return  455 ;
      when  473  => return  456 ;
      when  474  => return  456 ;
      when  475  => return  457 ;
      when  476  => return  458 ;
      when  477  => return  459 ;
      when  478  => return  460 ;
      when  479  => return  461 ;
      when  480  => return  462 ;
      when  481  => return  463 ;
      when  482  => return  464 ;
      when  483  => return  464 ;
      when  484  => return  465 ;
      when  485  => return  466 ;
      when  486  => return  467 ;
      when  487  => return  468 ;
      when  488  => return  469 ;
      when  489  => return  470 ;
      when  490  => return  471 ;
      when  491  => return  472 ;
      when  492  => return  472 ;
      when  493  => return  473 ;
      when  494  => return  474 ;
      when  495  => return  475 ;
      when  496  => return  476 ;
      when  497  => return  477 ;
      when  498  => return  478 ;
      when  499  => return  479 ;
      when  500  => return  479 ;
      when  501  => return  480 ;
      when  502  => return  481 ;
      when  503  => return  482 ;
      when  504  => return  483 ;
      when  505  => return  484 ;
      when  506  => return  485 ;
      when  507  => return  486 ;
      when  508  => return  486 ;
      when  509  => return  487 ;
      when  510  => return  488 ;
      when  511  => return  489 ;
      when  512  => return  490 ;
      when  513  => return  491 ;
      when  514  => return  492 ;
      when  515  => return  493 ;
      when  516  => return  493 ;
      when  517  => return  494 ;
      when  518  => return  495 ;
      when  519  => return  496 ;
      when  520  => return  497 ;
      when  521  => return  498 ;
      when  522  => return  499 ;
      when  523  => return  499 ;
      when  524  => return  500 ;
      when  525  => return  501 ;
      when  526  => return  502 ;
      when  527  => return  503 ;
      when  528  => return  504 ;
      when  529  => return  505 ;
      when  530  => return  506 ;
      when  531  => return  506 ;
      when  532  => return  507 ;
      when  533  => return  508 ;
      when  534  => return  509 ;
      when  535  => return  510 ;
      when  536  => return  511 ;
      when  537  => return  512 ;
      when  538  => return  512 ;
      when  539  => return  513 ;
      when  540  => return  514 ;
      when  541  => return  515 ;
      when  542  => return  516 ;
      when  543  => return  517 ;
      when  544  => return  518 ;
      when  545  => return  518 ;
      when  546  => return  519 ;
      when  547  => return  520 ;
      when  548  => return  521 ;
      when  549  => return  522 ;
      when  550  => return  523 ;
      when  551  => return  524 ;
      when  552  => return  524 ;
      when  553  => return  525 ;
      when  554  => return  526 ;
      when  555  => return  527 ;
      when  556  => return  528 ;
      when  557  => return  529 ;
      when  558  => return  529 ;
      when  559  => return  530 ;
      when  560  => return  531 ;
      when  561  => return  532 ;
      when  562  => return  533 ;
      when  563  => return  534 ;
      when  564  => return  535 ;
      when  565  => return  535 ;
      when  566  => return  536 ;
      when  567  => return  537 ;
      when  568  => return  538 ;
      when  569  => return  539 ;
      when  570  => return  540 ;
      when  571  => return  540 ;
      when  572  => return  541 ;
      when  573  => return  542 ;
      when  574  => return  543 ;
      when  575  => return  544 ;
      when  576  => return  545 ;
      when  577  => return  546 ;
      when  578  => return  546 ;
      when  579  => return  547 ;
      when  580  => return  548 ;
      when  581  => return  549 ;
      when  582  => return  550 ;
      when  583  => return  551 ;
      when  584  => return  551 ;
      when  585  => return  552 ;
      when  586  => return  553 ;
      when  587  => return  554 ;
      when  588  => return  555 ;
      when  589  => return  556 ;
      when  590  => return  556 ;
      when  591  => return  557 ;
      when  592  => return  558 ;
      when  593  => return  559 ;
      when  594  => return  560 ;
      when  595  => return  561 ;
      when  596  => return  561 ;
      when  597  => return  562 ;
      when  598  => return  563 ;
      when  599  => return  564 ;
      when  600  => return  565 ;
      when  601  => return  565 ;
      when  602  => return  566 ;
      when  603  => return  567 ;
      when  604  => return  568 ;
      when  605  => return  569 ;
      when  606  => return  570 ;
      when  607  => return  570 ;
      when  608  => return  571 ;
      when  609  => return  572 ;
      when  610  => return  573 ;
      when  611  => return  574 ;
      when  612  => return  575 ;
      when  613  => return  575 ;
      when  614  => return  576 ;
      when  615  => return  577 ;
      when  616  => return  578 ;
      when  617  => return  579 ;
      when  618  => return  579 ;
      when  619  => return  580 ;
      when  620  => return  581 ;
      when  621  => return  582 ;
      when  622  => return  583 ;
      when  623  => return  583 ;
      when  624  => return  584 ;
      when  625  => return  585 ;
      when  626  => return  586 ;
      when  627  => return  587 ;
      when  628  => return  588 ;
      when  629  => return  588 ;
      when  630  => return  589 ;
      when  631  => return  590 ;
      when  632  => return  591 ;
      when  633  => return  592 ;
      when  634  => return  592 ;
      when  635  => return  593 ;
      when  636  => return  594 ;
      when  637  => return  595 ;
      when  638  => return  596 ;
      when  639  => return  596 ;
      when  640  => return  597 ;
      when  641  => return  598 ;
      when  642  => return  599 ;
      when  643  => return  600 ;
      when  644  => return  600 ;
      when  645  => return  601 ;
      when  646  => return  602 ;
      when  647  => return  603 ;
      when  648  => return  604 ;
      when  649  => return  604 ;
      when  650  => return  605 ;
      when  651  => return  606 ;
      when  652  => return  607 ;
      when  653  => return  608 ;
      when  654  => return  608 ;
      when  655  => return  609 ;
      when  656  => return  610 ;
      when  657  => return  611 ;
      when  658  => return  612 ;
      when  659  => return  612 ;
      when  660  => return  613 ;
      when  661  => return  614 ;
      when  662  => return  615 ;
      when  663  => return  615 ;
      when  664  => return  616 ;
      when  665  => return  617 ;
      when  666  => return  618 ;
      when  667  => return  619 ;
      when  668  => return  619 ;
      when  669  => return  620 ;
      when  670  => return  621 ;
      when  671  => return  622 ;
      when  672  => return  623 ;
      when  673  => return  623 ;
      when  674  => return  624 ;
      when  675  => return  625 ;
      when  676  => return  626 ;
      when  677  => return  626 ;
      when  678  => return  627 ;
      when  679  => return  628 ;
      when  680  => return  629 ;
      when  681  => return  630 ;
      when  682  => return  630 ;
      when  683  => return  631 ;
      when  684  => return  632 ;
      when  685  => return  633 ;
      when  686  => return  633 ;
      when  687  => return  634 ;
      when  688  => return  635 ;
      when  689  => return  636 ;
      when  690  => return  637 ;
      when  691  => return  637 ;
      when  692  => return  638 ;
      when  693  => return  639 ;
      when  694  => return  640 ;
      when  695  => return  640 ;
      when  696  => return  641 ;
      when  697  => return  642 ;
      when  698  => return  643 ;
      when  699  => return  643 ;
      when  700  => return  644 ;
      when  701  => return  645 ;
      when  702  => return  646 ;
      when  703  => return  647 ;
      when  704  => return  647 ;
      when  705  => return  648 ;
      when  706  => return  649 ;
      when  707  => return  650 ;
      when  708  => return  650 ;
      when  709  => return  651 ;
      when  710  => return  652 ;
      when  711  => return  653 ;
      when  712  => return  653 ;
      when  713  => return  654 ;
      when  714  => return  655 ;
      when  715  => return  656 ;
      when  716  => return  656 ;
      when  717  => return  657 ;
      when  718  => return  658 ;
      when  719  => return  659 ;
      when  720  => return  659 ;
      when  721  => return  660 ;
      when  722  => return  661 ;
      when  723  => return  662 ;
      when  724  => return  662 ;
      when  725  => return  663 ;
      when  726  => return  664 ;
      when  727  => return  665 ;
      when  728  => return  665 ;
      when  729  => return  666 ;
      when  730  => return  667 ;
      when  731  => return  668 ;
      when  732  => return  668 ;
      when  733  => return  669 ;
      when  734  => return  670 ;
      when  735  => return  671 ;
      when  736  => return  671 ;
      when  737  => return  672 ;
      when  738  => return  673 ;
      when  739  => return  674 ;
      when  740  => return  674 ;
      when  741  => return  675 ;
      when  742  => return  676 ;
      when  743  => return  677 ;
      when  744  => return  677 ;
      when  745  => return  678 ;
      when  746  => return  679 ;
      when  747  => return  679 ;
      when  748  => return  680 ;
      when  749  => return  681 ;
      when  750  => return  682 ;
      when  751  => return  682 ;
      when  752  => return  683 ;
      when  753  => return  684 ;
      when  754  => return  685 ;
      when  755  => return  685 ;
      when  756  => return  686 ;
      when  757  => return  687 ;
      when  758  => return  687 ;
      when  759  => return  688 ;
      when  760  => return  689 ;
      when  761  => return  690 ;
      when  762  => return  690 ;
      when  763  => return  691 ;
      when  764  => return  692 ;
      when  765  => return  693 ;
      when  766  => return  693 ;
      when  767  => return  694 ;
      when  768  => return  695 ;
      when  769  => return  695 ;
      when  770  => return  696 ;
      when  771  => return  697 ;
      when  772  => return  698 ;
      when  773  => return  698 ;
      when  774  => return  699 ;
      when  775  => return  700 ;
      when  776  => return  700 ;
      when  777  => return  701 ;
      when  778  => return  702 ;
      when  779  => return  703 ;
      when  780  => return  703 ;
      when  781  => return  704 ;
      when  782  => return  705 ;
      when  783  => return  705 ;
      when  784  => return  706 ;
      when  785  => return  707 ;
      when  786  => return  708 ;
      when  787  => return  708 ;
      when  788  => return  709 ;
      when  789  => return  710 ;
      when  790  => return  710 ;
      when  791  => return  711 ;
      when  792  => return  712 ;
      when  793  => return  712 ;
      when  794  => return  713 ;
      when  795  => return  714 ;
      when  796  => return  715 ;
      when  797  => return  715 ;
      when  798  => return  716 ;
      when  799  => return  717 ;
      when  800  => return  717 ;
      when  801  => return  718 ;
      when  802  => return  719 ;
      when  803  => return  719 ;
      when  804  => return  720 ;
      when  805  => return  721 ;
      when  806  => return  722 ;
      when  807  => return  722 ;
      when  808  => return  723 ;
      when  809  => return  724 ;
      when  810  => return  724 ;
      when  811  => return  725 ;
      when  812  => return  726 ;
      when  813  => return  726 ;
      when  814  => return  727 ;
      when  815  => return  728 ;
      when  816  => return  728 ;
      when  817  => return  729 ;
      when  818  => return  730 ;
      when  819  => return  730 ;
      when  820  => return  731 ;
      when  821  => return  732 ;
      when  822  => return  733 ;
      when  823  => return  733 ;
      when  824  => return  734 ;
      when  825  => return  735 ;
      when  826  => return  735 ;
      when  827  => return  736 ;
      when  828  => return  737 ;
      when  829  => return  737 ;
      when  830  => return  738 ;
      when  831  => return  739 ;
      when  832  => return  739 ;
      when  833  => return  740 ;
      when  834  => return  741 ;
      when  835  => return  741 ;
      when  836  => return  742 ;
      when  837  => return  743 ;
      when  838  => return  743 ;
      when  839  => return  744 ;
      when  840  => return  745 ;
      when  841  => return  745 ;
      when  842  => return  746 ;
      when  843  => return  747 ;
      when  844  => return  747 ;
      when  845  => return  748 ;
      when  846  => return  749 ;
      when  847  => return  749 ;
      when  848  => return  750 ;
      when  849  => return  751 ;
      when  850  => return  751 ;
      when  851  => return  752 ;
      when  852  => return  753 ;
      when  853  => return  753 ;
      when  854  => return  754 ;
      when  855  => return  755 ;
      when  856  => return  755 ;
      when  857  => return  756 ;
      when  858  => return  757 ;
      when  859  => return  757 ;
      when  860  => return  758 ;
      when  861  => return  758 ;
      when  862  => return  759 ;
      when  863  => return  760 ;
      when  864  => return  760 ;
      when  865  => return  761 ;
      when  866  => return  762 ;
      when  867  => return  762 ;
      when  868  => return  763 ;
      when  869  => return  764 ;
      when  870  => return  764 ;
      when  871  => return  765 ;
      when  872  => return  766 ;
      when  873  => return  766 ;
      when  874  => return  767 ;
      when  875  => return  768 ;
      when  876  => return  768 ;
      when  877  => return  769 ;
      when  878  => return  769 ;
      when  879  => return  770 ;
      when  880  => return  771 ;
      when  881  => return  771 ;
      when  882  => return  772 ;
      when  883  => return  773 ;
      when  884  => return  773 ;
      when  885  => return  774 ;
      when  886  => return  775 ;
      when  887  => return  775 ;
      when  888  => return  776 ;
      when  889  => return  776 ;
      when  890  => return  777 ;
      when  891  => return  778 ;
      when  892  => return  778 ;
      when  893  => return  779 ;
      when  894  => return  780 ;
      when  895  => return  780 ;
      when  896  => return  781 ;
      when  897  => return  781 ;
      when  898  => return  782 ;
      when  899  => return  783 ;
      when  900  => return  783 ;
      when  901  => return  784 ;
      when  902  => return  785 ;
      when  903  => return  785 ;
      when  904  => return  786 ;
      when  905  => return  786 ;
      when  906  => return  787 ;
      when  907  => return  788 ;
      when  908  => return  788 ;
      when  909  => return  789 ;
      when  910  => return  790 ;
      when  911  => return  790 ;
      when  912  => return  791 ;
      when  913  => return  791 ;
      when  914  => return  792 ;
      when  915  => return  793 ;
      when  916  => return  793 ;
      when  917  => return  794 ;
      when  918  => return  794 ;
      when  919  => return  795 ;
      when  920  => return  796 ;
      when  921  => return  796 ;
      when  922  => return  797 ;
      when  923  => return  797 ;
      when  924  => return  798 ;
      when  925  => return  799 ;
      when  926  => return  799 ;
      when  927  => return  800 ;
      when  928  => return  800 ;
      when  929  => return  801 ;
      when  930  => return  802 ;
      when  931  => return  802 ;
      when  932  => return  803 ;
      when  933  => return  803 ;
      when  934  => return  804 ;
      when  935  => return  805 ;
      when  936  => return  805 ;
      when  937  => return  806 ;
      when  938  => return  806 ;
      when  939  => return  807 ;
      when  940  => return  808 ;
      when  941  => return  808 ;
      when  942  => return  809 ;
      when  943  => return  809 ;
      when  944  => return  810 ;
      when  945  => return  810 ;
      when  946  => return  811 ;
      when  947  => return  812 ;
      when  948  => return  812 ;
      when  949  => return  813 ;
      when  950  => return  813 ;
      when  951  => return  814 ;
      when  952  => return  815 ;
      when  953  => return  815 ;
      when  954  => return  816 ;
      when  955  => return  816 ;
      when  956  => return  817 ;
      when  957  => return  817 ;
      when  958  => return  818 ;
      when  959  => return  819 ;
      when  960  => return  819 ;
      when  961  => return  820 ;
      when  962  => return  820 ;
      when  963  => return  821 ;
      when  964  => return  821 ;
      when  965  => return  822 ;
      when  966  => return  823 ;
      when  967  => return  823 ;
      when  968  => return  824 ;
      when  969  => return  824 ;
      when  970  => return  825 ;
      when  971  => return  825 ;
      when  972  => return  826 ;
      when  973  => return  827 ;
      when  974  => return  827 ;
      when  975  => return  828 ;
      when  976  => return  828 ;
      when  977  => return  829 ;
      when  978  => return  829 ;
      when  979  => return  830 ;
      when  980  => return  830 ;
      when  981  => return  831 ;
      when  982  => return  832 ;
      when  983  => return  832 ;
      when  984  => return  833 ;
      when  985  => return  833 ;
      when  986  => return  834 ;
      when  987  => return  834 ;
      when  988  => return  835 ;
      when  989  => return  835 ;
      when  990  => return  836 ;
      when  991  => return  837 ;
      when  992  => return  837 ;
      when  993  => return  838 ;
      when  994  => return  838 ;
      when  995  => return  839 ;
      when  996  => return  839 ;
      when  997  => return  840 ;
      when  998  => return  840 ;
      when  999  => return  841 ;
      when  1000  => return  841 ;
      when  1001  => return  842 ;
      when  1002  => return  843 ;
      when  1003  => return  843 ;
      when  1004  => return  844 ;
      when  1005  => return  844 ;
      when  1006  => return  845 ;
      when  1007  => return  845 ;
      when  1008  => return  846 ;
      when  1009  => return  846 ;
      when  1010  => return  847 ;
      when  1011  => return  847 ;
      when  1012  => return  848 ;
      when  1013  => return  848 ;
      when  1014  => return  849 ;
      when  1015  => return  849 ;
      when  1016  => return  850 ;
      when  1017  => return  851 ;
      when  1018  => return  851 ;
      when  1019  => return  852 ;
      when  1020  => return  852 ;
      when  1021  => return  853 ;
      when  1022  => return  853 ;
      when  1023  => return  854 ;
      when  1024  => return  854 ;
      when  1025  => return  855 ;
      when  1026  => return  855 ;
      when  1027  => return  856 ;
      when  1028  => return  856 ;
      when  1029  => return  857 ;
      when  1030  => return  857 ;
      when  1031  => return  858 ;
      when  1032  => return  858 ;
      when  1033  => return  859 ;
      when  1034  => return  859 ;
      when  1035  => return  860 ;
      when  1036  => return  860 ;
      when  1037  => return  861 ;
      when  1038  => return  861 ;
      when  1039  => return  862 ;
      when  1040  => return  862 ;
      when  1041  => return  863 ;
      when  1042  => return  863 ;
      when  1043  => return  864 ;
      when  1044  => return  864 ;
      when  1045  => return  865 ;
      when  1046  => return  865 ;
      when  1047  => return  866 ;
      when  1048  => return  866 ;
      when  1049  => return  867 ;
      when  1050  => return  867 ;
      when  1051  => return  868 ;
      when  1052  => return  868 ;
      when  1053  => return  869 ;
      when  1054  => return  869 ;
      when  1055  => return  870 ;
      when  1056  => return  870 ;
      when  1057  => return  871 ;
      when  1058  => return  871 ;
      when  1059  => return  872 ;
      when  1060  => return  872 ;
      when  1061  => return  873 ;
      when  1062  => return  873 ;
      when  1063  => return  874 ;
      when  1064  => return  874 ;
      when  1065  => return  875 ;
      when  1066  => return  875 ;
      when  1067  => return  876 ;
      when  1068  => return  876 ;
      when  1069  => return  877 ;
      when  1070  => return  877 ;
      when  1071  => return  878 ;
      when  1072  => return  878 ;
      when  1073  => return  879 ;
      when  1074  => return  879 ;
      when  1075  => return  880 ;
      when  1076  => return  880 ;
      when  1077  => return  881 ;
      when  1078  => return  881 ;
      when  1079  => return  881 ;
      when  1080  => return  882 ;
      when  1081  => return  882 ;
      when  1082  => return  883 ;
      when  1083  => return  883 ;
      when  1084  => return  884 ;
      when  1085  => return  884 ;
      when  1086  => return  885 ;
      when  1087  => return  885 ;
      when  1088  => return  886 ;
      when  1089  => return  886 ;
      when  1090  => return  887 ;
      when  1091  => return  887 ;
      when  1092  => return  888 ;
      when  1093  => return  888 ;
      when  1094  => return  888 ;
      when  1095  => return  889 ;
      when  1096  => return  889 ;
      when  1097  => return  890 ;
      when  1098  => return  890 ;
      when  1099  => return  891 ;
      when  1100  => return  891 ;
      when  1101  => return  892 ;
      when  1102  => return  892 ;
      when  1103  => return  893 ;
      when  1104  => return  893 ;
      when  1105  => return  893 ;
      when  1106  => return  894 ;
      when  1107  => return  894 ;
      when  1108  => return  895 ;
      when  1109  => return  895 ;
      when  1110  => return  896 ;
      when  1111  => return  896 ;
      when  1112  => return  897 ;
      when  1113  => return  897 ;
      when  1114  => return  897 ;
      when  1115  => return  898 ;
      when  1116  => return  898 ;
      when  1117  => return  899 ;
      when  1118  => return  899 ;
      when  1119  => return  900 ;
      when  1120  => return  900 ;
      when  1121  => return  901 ;
      when  1122  => return  901 ;
      when  1123  => return  901 ;
      when  1124  => return  902 ;
      when  1125  => return  902 ;
      when  1126  => return  903 ;
      when  1127  => return  903 ;
      when  1128  => return  904 ;
      when  1129  => return  904 ;
      when  1130  => return  904 ;
      when  1131  => return  905 ;
      when  1132  => return  905 ;
      when  1133  => return  906 ;
      when  1134  => return  906 ;
      when  1135  => return  907 ;
      when  1136  => return  907 ;
      when  1137  => return  907 ;
      when  1138  => return  908 ;
      when  1139  => return  908 ;
      when  1140  => return  909 ;
      when  1141  => return  909 ;
      when  1142  => return  909 ;
      when  1143  => return  910 ;
      when  1144  => return  910 ;
      when  1145  => return  911 ;
      when  1146  => return  911 ;
      when  1147  => return  912 ;
      when  1148  => return  912 ;
      when  1149  => return  912 ;
      when  1150  => return  913 ;
      when  1151  => return  913 ;
      when  1152  => return  914 ;
      when  1153  => return  914 ;
      when  1154  => return  914 ;
      when  1155  => return  915 ;
      when  1156  => return  915 ;
      when  1157  => return  916 ;
      when  1158  => return  916 ;
      when  1159  => return  916 ;
      when  1160  => return  917 ;
      when  1161  => return  917 ;
      when  1162  => return  918 ;
      when  1163  => return  918 ;
      when  1164  => return  918 ;
      when  1165  => return  919 ;
      when  1166  => return  919 ;
      when  1167  => return  920 ;
      when  1168  => return  920 ;
      when  1169  => return  920 ;
      when  1170  => return  921 ;
      when  1171  => return  921 ;
      when  1172  => return  922 ;
      when  1173  => return  922 ;
      when  1174  => return  922 ;
      when  1175  => return  923 ;
      when  1176  => return  923 ;
      when  1177  => return  923 ;
      when  1178  => return  924 ;
      when  1179  => return  924 ;
      when  1180  => return  925 ;
      when  1181  => return  925 ;
      when  1182  => return  925 ;
      when  1183  => return  926 ;
      when  1184  => return  926 ;
      when  1185  => return  926 ;
      when  1186  => return  927 ;
      when  1187  => return  927 ;
      when  1188  => return  928 ;
      when  1189  => return  928 ;
      when  1190  => return  928 ;
      when  1191  => return  929 ;
      when  1192  => return  929 ;
      when  1193  => return  929 ;
      when  1194  => return  930 ;
      when  1195  => return  930 ;
      when  1196  => return  931 ;
      when  1197  => return  931 ;
      when  1198  => return  931 ;
      when  1199  => return  932 ;
      when  1200  => return  932 ;
      when  1201  => return  932 ;
      when  1202  => return  933 ;
      when  1203  => return  933 ;
      when  1204  => return  933 ;
      when  1205  => return  934 ;
      when  1206  => return  934 ;
      when  1207  => return  935 ;
      when  1208  => return  935 ;
      when  1209  => return  935 ;
      when  1210  => return  936 ;
      when  1211  => return  936 ;
      when  1212  => return  936 ;
      when  1213  => return  937 ;
      when  1214  => return  937 ;
      when  1215  => return  937 ;
      when  1216  => return  938 ;
      when  1217  => return  938 ;
      when  1218  => return  938 ;
      when  1219  => return  939 ;
      when  1220  => return  939 ;
      when  1221  => return  939 ;
      when  1222  => return  940 ;
      when  1223  => return  940 ;
      when  1224  => return  940 ;
      when  1225  => return  941 ;
      when  1226  => return  941 ;
      when  1227  => return  941 ;
      when  1228  => return  942 ;
      when  1229  => return  942 ;
      when  1230  => return  942 ;
      when  1231  => return  943 ;
      when  1232  => return  943 ;
      when  1233  => return  943 ;
      when  1234  => return  944 ;
      when  1235  => return  944 ;
      when  1236  => return  944 ;
      when  1237  => return  945 ;
      when  1238  => return  945 ;
      when  1239  => return  945 ;
      when  1240  => return  946 ;
      when  1241  => return  946 ;
      when  1242  => return  946 ;
      when  1243  => return  947 ;
      when  1244  => return  947 ;
      when  1245  => return  947 ;
      when  1246  => return  948 ;
      when  1247  => return  948 ;
      when  1248  => return  948 ;
      when  1249  => return  949 ;
      when  1250  => return  949 ;
      when  1251  => return  949 ;
      when  1252  => return  950 ;
      when  1253  => return  950 ;
      when  1254  => return  950 ;
      when  1255  => return  951 ;
      when  1256  => return  951 ;
      when  1257  => return  951 ;
      when  1258  => return  951 ;
      when  1259  => return  952 ;
      when  1260  => return  952 ;
      when  1261  => return  952 ;
      when  1262  => return  953 ;
      when  1263  => return  953 ;
      when  1264  => return  953 ;
      when  1265  => return  954 ;
      when  1266  => return  954 ;
      when  1267  => return  954 ;
      when  1268  => return  955 ;
      when  1269  => return  955 ;
      when  1270  => return  955 ;
      when  1271  => return  955 ;
      when  1272  => return  956 ;
      when  1273  => return  956 ;
      when  1274  => return  956 ;
      when  1275  => return  957 ;
      when  1276  => return  957 ;
      when  1277  => return  957 ;
      when  1278  => return  957 ;
      when  1279  => return  958 ;
      when  1280  => return  958 ;
      when  1281  => return  958 ;
      when  1282  => return  959 ;
      when  1283  => return  959 ;
      when  1284  => return  959 ;
      when  1285  => return  959 ;
      when  1286  => return  960 ;
      when  1287  => return  960 ;
      when  1288  => return  960 ;
      when  1289  => return  961 ;
      when  1290  => return  961 ;
      when  1291  => return  961 ;
      when  1292  => return  961 ;
      when  1293  => return  962 ;
      when  1294  => return  962 ;
      when  1295  => return  962 ;
      when  1296  => return  962 ;
      when  1297  => return  963 ;
      when  1298  => return  963 ;
      when  1299  => return  963 ;
      when  1300  => return  964 ;
      when  1301  => return  964 ;
      when  1302  => return  964 ;
      when  1303  => return  964 ;
      when  1304  => return  965 ;
      when  1305  => return  965 ;
      when  1306  => return  965 ;
      when  1307  => return  965 ;
      when  1308  => return  966 ;
      when  1309  => return  966 ;
      when  1310  => return  966 ;
      when  1311  => return  966 ;
      when  1312  => return  967 ;
      when  1313  => return  967 ;
      when  1314  => return  967 ;
      when  1315  => return  967 ;
      when  1316  => return  968 ;
      when  1317  => return  968 ;
      when  1318  => return  968 ;
      when  1319  => return  968 ;
      when  1320  => return  969 ;
      when  1321  => return  969 ;
      when  1322  => return  969 ;
      when  1323  => return  969 ;
      when  1324  => return  970 ;
      when  1325  => return  970 ;
      when  1326  => return  970 ;
      when  1327  => return  970 ;
      when  1328  => return  971 ;
      when  1329  => return  971 ;
      when  1330  => return  971 ;
      when  1331  => return  971 ;
      when  1332  => return  972 ;
      when  1333  => return  972 ;
      when  1334  => return  972 ;
      when  1335  => return  972 ;
      when  1336  => return  973 ;
      when  1337  => return  973 ;
      when  1338  => return  973 ;
      when  1339  => return  973 ;
      when  1340  => return  973 ;
      when  1341  => return  974 ;
      when  1342  => return  974 ;
      when  1343  => return  974 ;
      when  1344  => return  974 ;
      when  1345  => return  975 ;
      when  1346  => return  975 ;
      when  1347  => return  975 ;
      when  1348  => return  975 ;
      when  1349  => return  976 ;
      when  1350  => return  976 ;
      when  1351  => return  976 ;
      when  1352  => return  976 ;
      when  1353  => return  976 ;
      when  1354  => return  977 ;
      when  1355  => return  977 ;
      when  1356  => return  977 ;
      when  1357  => return  977 ;
      when  1358  => return  977 ;
      when  1359  => return  978 ;
      when  1360  => return  978 ;
      when  1361  => return  978 ;
      when  1362  => return  978 ;
      when  1363  => return  978 ;
      when  1364  => return  979 ;
      when  1365  => return  979 ;
      when  1366  => return  979 ;
      when  1367  => return  979 ;
      when  1368  => return  980 ;
      when  1369  => return  980 ;
      when  1370  => return  980 ;
      when  1371  => return  980 ;
      when  1372  => return  980 ;
      when  1373  => return  981 ;
      when  1374  => return  981 ;
      when  1375  => return  981 ;
      when  1376  => return  981 ;
      when  1377  => return  981 ;
      when  1378  => return  981 ;
      when  1379  => return  982 ;
      when  1380  => return  982 ;
      when  1381  => return  982 ;
      when  1382  => return  982 ;
      when  1383  => return  982 ;
      when  1384  => return  983 ;
      when  1385  => return  983 ;
      when  1386  => return  983 ;
      when  1387  => return  983 ;
      when  1388  => return  983 ;
      when  1389  => return  984 ;
      when  1390  => return  984 ;
      when  1391  => return  984 ;
      when  1392  => return  984 ;
      when  1393  => return  984 ;
      when  1394  => return  984 ;
      when  1395  => return  985 ;
      when  1396  => return  985 ;
      when  1397  => return  985 ;
      when  1398  => return  985 ;
      when  1399  => return  985 ;
      when  1400  => return  985 ;
      when  1401  => return  986 ;
      when  1402  => return  986 ;
      when  1403  => return  986 ;
      when  1404  => return  986 ;
      when  1405  => return  986 ;
      when  1406  => return  986 ;
      when  1407  => return  987 ;
      when  1408  => return  987 ;
      when  1409  => return  987 ;
      when  1410  => return  987 ;
      when  1411  => return  987 ;
      when  1412  => return  987 ;
      when  1413  => return  988 ;
      when  1414  => return  988 ;
      when  1415  => return  988 ;
      when  1416  => return  988 ;
      when  1417  => return  988 ;
      when  1418  => return  988 ;
      when  1419  => return  989 ;
      when  1420  => return  989 ;
      when  1421  => return  989 ;
      when  1422  => return  989 ;
      when  1423  => return  989 ;
      when  1424  => return  989 ;
      when  1425  => return  989 ;
      when  1426  => return  990 ;
      when  1427  => return  990 ;
      when  1428  => return  990 ;
      when  1429  => return  990 ;
      when  1430  => return  990 ;
      when  1431  => return  990 ;
      when  1432  => return  990 ;
      when  1433  => return  991 ;
      when  1434  => return  991 ;
      when  1435  => return  991 ;
      when  1436  => return  991 ;
      when  1437  => return  991 ;
      when  1438  => return  991 ;
      when  1439  => return  991 ;
      when  1440  => return  991 ;
      when  1441  => return  992 ;
      when  1442  => return  992 ;
      when  1443  => return  992 ;
      when  1444  => return  992 ;
      when  1445  => return  992 ;
      when  1446  => return  992 ;
      when  1447  => return  992 ;
      when  1448  => return  992 ;
      when  1449  => return  993 ;
      when  1450  => return  993 ;
      when  1451  => return  993 ;
      when  1452  => return  993 ;
      when  1453  => return  993 ;
      when  1454  => return  993 ;
      when  1455  => return  993 ;
      when  1456  => return  993 ;
      when  1457  => return  994 ;
      when  1458  => return  994 ;
      when  1459  => return  994 ;
      when  1460  => return  994 ;
      when  1461  => return  994 ;
      when  1462  => return  994 ;
      when  1463  => return  994 ;
      when  1464  => return  994 ;
      when  1465  => return  994 ;
      when  1466  => return  995 ;
      when  1467  => return  995 ;
      when  1468  => return  995 ;
      when  1469  => return  995 ;
      when  1470  => return  995 ;
      when  1471  => return  995 ;
      when  1472  => return  995 ;
      when  1473  => return  995 ;
      when  1474  => return  995 ;
      when  1475  => return  995 ;
      when  1476  => return  996 ;
      when  1477  => return  996 ;
      when  1478  => return  996 ;
      when  1479  => return  996 ;
      when  1480  => return  996 ;
      when  1481  => return  996 ;
      when  1482  => return  996 ;
      when  1483  => return  996 ;
      when  1484  => return  996 ;
      when  1485  => return  996 ;
      when  1486  => return  996 ;
      when  1487  => return  996 ;
      when  1488  => return  997 ;
      when  1489  => return  997 ;
      when  1490  => return  997 ;
      when  1491  => return  997 ;
      when  1492  => return  997 ;
      when  1493  => return  997 ;
      when  1494  => return  997 ;
      when  1495  => return  997 ;
      when  1496  => return  997 ;
      when  1497  => return  997 ;
      when  1498  => return  997 ;
      when  1499  => return  997 ;
      when  1500  => return  997 ;
      when  1501  => return  998 ;
      when  1502  => return  998 ;
      when  1503  => return  998 ;
      when  1504  => return  998 ;
      when  1505  => return  998 ;
      when  1506  => return  998 ;
      when  1507  => return  998 ;
      when  1508  => return  998 ;
      when  1509  => return  998 ;
      when  1510  => return  998 ;
      when  1511  => return  998 ;
      when  1512  => return  998 ;
      when  1513  => return  998 ;
      when  1514  => return  998 ;
      when  1515  => return  998 ;
      when  1516  => return  998 ;
      when  1517  => return  999 ;
      when  1518  => return  999 ;
      when  1519  => return  999 ;
      when  1520  => return  999 ;
      when  1521  => return  999 ;
      when  1522  => return  999 ;
      when  1523  => return  999 ;
      when  1524  => return  999 ;
      when  1525  => return  999 ;
      when  1526  => return  999 ;
      when  1527  => return  999 ;
      when  1528  => return  999 ;
      when  1529  => return  999 ;
      when  1530  => return  999 ;
      when  1531  => return  999 ;
      when  1532  => return  999 ;
      when  1533  => return  999 ;
      when  1534  => return  999 ;
      when  1535  => return  999 ;
      when  1536  => return  999 ;
      when  1537  => return  999 ;
      when  1538  => return  999 ;
      when  1539  => return  999 ;
      when  1540  => return  1000 ;
      when  1541  => return  1000 ;
      when  1542  => return  1000 ;
      when  1543  => return  1000 ;
      when  1544  => return  1000 ;
      when  1545  => return  1000 ;
      when  1546  => return  1000 ;
      when  1547  => return  1000 ;
      when  1548  => return  1000 ;
      when  1549  => return  1000 ;
      when  1550  => return  1000 ;
      when  1551  => return  1000 ;
      when  1552  => return  1000 ;
      when  1553  => return  1000 ;
      when  1554  => return  1000 ;
      when  1555  => return  1000 ;
      when  1556  => return  1000 ;
      when  1557  => return  1000 ;
      when  1558  => return  1000 ;
      when  1559  => return  1000 ;
      when  1560  => return  1000 ;
      when  1561  => return  1000 ;
      when  1562  => return  1000 ;
      when  1563  => return  1000 ;
      when  1564  => return  1000 ;
      when  1565  => return  1000 ;
      when  1566  => return  1000 ;
      when  1567  => return  1000 ;
      when  1568  => return  1000 ;
      when  1569  => return  1000 ;
		when others => return 0;
    end case;
  end function;

  function sin(x : integer ) return integer is
  begin
    case div(x, pi/2) is
      when 0 =>
        return sin_0_pi2(x);
      when 1 =>
        return sin_0_pi2(x-pi);
      when 2 =>
        return -1*sin_0_pi2(x);
      when others =>
        return -1*sin_0_pi2(x-pi); --depois checar se nao ocorre underflow aqui
    end case;
  end function;

begin
  increment_t: process(clk)
  begin
    if rising_edge(clk) then
      t := (t + 1);
		x_tmp := std_logic_vector(to_signed(x_ampl * sin(t + alpha + delta),16));
		y_tmp := std_logic_vector(to_signed(y_ampl * sin(t + beta),16));
    end if;
  end process;

  x_out <= x_tmp;
  y_out <= y_tmp;
end arq;
